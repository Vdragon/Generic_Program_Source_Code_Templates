// 〈程式檔名〉 - 〈程式描述文字（一言以蔽之）〉
// 〈程式智慧財產權擁有者名諱、地址（選用）〉 © 〈智慧財產權生效年〉

//時脈產生器半週期
//`define CLOCK_PERIOD_HALF 10

module module_name();
//宣告port類型
  output reg ;
  input wire ;

	//D.U.T. instantiation

  /* 時脈產生器
  always begin
    #`CLOCK_PERIOD_HALF Clk = !Clk;
	end
  */
  
  initial begin

	end
endmodule